library IEEE;
use IEEE.STD_LOGIC_1164.all;

package trc_packages is
  -- Define your 2D array type here
  type vector_of_vectors is array (natural range <>) of std_logic_vector;
end package trc_packages;
